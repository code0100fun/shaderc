module shaderc
