module shaderc

#flag -L @VMODROOT/thirdparty/build/shaderc/libshaderc/
#flag -I @VMODROOT/thirdparty/shaderc/libshaderc/include
#flag -llibshaderc_shared
#include "shaderc/shaderc.h"
