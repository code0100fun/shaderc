module shaderc

#flag -L @VMODROOT/build/shaderc/libshaderc
#flag -I @VMODROOT/thirdparty/shaderc/libshaderc/include
#flag -lshaderc_shared
#include "shaderc/shaderc.h"
